`define RST1_CYCLE_NUM 10
`define RST0_CYCLE_NUM 60