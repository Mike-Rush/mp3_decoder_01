`define RST_CYCLE_NUM 5